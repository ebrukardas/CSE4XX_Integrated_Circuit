magic
tech scmos
timestamp 1541705767
<< nwell >>
rect -44 -24 -16 -2
<< polysilicon >>
rect -36 -10 -34 -7
rect -26 -10 -24 -7
rect -36 -37 -34 -18
rect -26 -37 -24 -18
rect -36 -44 -34 -41
rect -26 -44 -24 -41
<< ndiffusion >>
rect -38 -41 -36 -37
rect -34 -41 -32 -37
rect -28 -41 -26 -37
rect -24 -41 -22 -37
<< pdiffusion >>
rect -38 -18 -36 -10
rect -34 -18 -26 -10
rect -24 -18 -22 -10
<< metal1 >>
rect -44 0 -16 1
rect -44 -4 -42 0
rect -38 -4 -16 0
rect -44 -5 -16 -4
rect -42 -10 -38 -5
rect -22 -22 -18 -18
rect -32 -26 -18 -22
rect -32 -37 -28 -26
rect -42 -46 -38 -41
rect -22 -46 -18 -41
rect -44 -47 -15 -46
rect -44 -51 -42 -47
rect -38 -51 -22 -47
rect -18 -51 -15 -47
rect -44 -52 -15 -51
<< ntransistor >>
rect -36 -41 -34 -37
rect -26 -41 -24 -37
<< ptransistor >>
rect -36 -18 -34 -10
rect -26 -18 -24 -10
<< polycontact >>
rect -40 -33 -36 -29
rect -24 -33 -20 -29
<< ndcontact >>
rect -42 -41 -38 -37
rect -32 -41 -28 -37
rect -22 -41 -18 -37
rect -42 -51 -38 -47
rect -22 -51 -18 -47
<< pdcontact >>
rect -42 -4 -38 0
rect -42 -18 -38 -10
rect -22 -18 -18 -10
<< labels >>
rlabel metal1 -30 0 -30 0 1 VDD
rlabel metal1 -19 -25 -19 -25 1 Vout
rlabel polycontact -38 -31 -38 -31 1 VinA
rlabel polycontact -22 -31 -22 -31 1 VinB
rlabel metal1 -31 -49 -31 -49 1 GND
<< end >>
