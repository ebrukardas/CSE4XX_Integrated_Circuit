* SPICE3 file created from mux_2.ext - technology: scmos

.option scale=0.12u

M1000 snot Vselk VDD w_n3_28# pmos w=8 l=2
+  ad=48 pd=28 as=320 ps=220
M1001 a_28_34# snot VDD w_n3_28# pmos w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1002 and1 Vin0 a_28_34# w_n3_28# pmos w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1003 GND and1 VDD w_n3_28# pmos w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1004 VDD and2 GND w_n3_28# pmos w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_84_34# Vin1 VDD w_n3_28# pmos w=8 l=2
+  ad=64 pd=32 as=0 ps=0
M1006 and2 Vselk a_84_34# w_n3_28# pmos w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1007 snot Vselk GND Gnd nmos w=4 l=2
+  ad=24 pd=20 as=264 ps=236
M1008 and1 snot GND Gnd nmos w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1009 GND Vin0 and1 Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_56_11# and1 GND Gnd nmos w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1011 GND and2 a_56_11# Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1012 and2 Vin1 GND Gnd nmos w=4 l=2
+  ad=32 pd=24 as=0 ps=0
M1013 GND Vselk and2 Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n3_28# and2 4.8fF
C1 w_n3_28# Vin0 2.6fF
C2 w_n3_28# Vselk 7.3fF
C3 w_n3_28# Vin1 2.6fF
C4 w_n3_28# VDD 16.6fF
C5 w_n3_28# snot 3.8fF
C6 and2 Vselk 0.2fF
C7 w_n3_28# and1 3.8fF
C8 and2 Vin1 0.2fF
C9 Vselk VDD 0.7fF
C10 Vin0 and1 0.2fF
C11 Vin1 Gnd 8.8fF
C12 and2 Gnd 11.1fF
C13 and1 Gnd 10.4fF
C14 Vin0 Gnd 8.8fF
C15 snot Gnd 9.1fF
C16 VDD Gnd 11.9fF
C17 Vselk Gnd 34.7fF
C18 w_n3_28# Gnd 1.1fF


*
* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    Vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2   V2   T3   V3   T4    V4    T5   V5    T5   V5     T5   V5     T5   V5 
*----- ----- ----- ------ --  --   ---  --   ---- --   ---   --    ---- --    ----  --    ----  --    ----  -- 
Vin0   Vin0   0    PWL(    0  0    3.9N  0   4N  2.5   7.9N  2.5   8N   0     11.9N  0     12N  2.5   15.9N  2.5  ) 
Vin1   Vin1   0    PWL(    0  0    3.9N  0   4N  0	   7.9N  0     8N   2.5   11.9N  2.5   12N  2.5   15.9N  2.5 )
Vselk   Vselk 0    PWL(    0  0    3.9N  0   4N  0	   7.9N  0     8N   2.5   11.9N  2.5   12N  2.5   15.9N  2.5 )


*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  20.2N


* The following line is for DC analysis

.DC VIN0 0 2.6 0.1

* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
