magic
tech scmos
timestamp 1542645901
<< nwell >>
rect -3 28 104 50
<< polysilicon >>
rect 5 57 94 59
rect 8 42 10 57
rect 26 42 28 45
rect 36 42 38 45
rect 54 42 56 45
rect 64 42 66 45
rect 82 42 84 45
rect 92 42 94 57
rect 8 15 10 34
rect 26 15 28 34
rect 36 15 38 34
rect 54 15 56 34
rect 64 15 66 34
rect 82 15 84 34
rect 92 15 94 34
rect 8 8 10 11
rect 26 8 28 11
rect 36 -3 38 11
rect 54 9 56 11
rect 64 9 66 11
rect 82 -3 84 11
rect 92 8 94 11
<< ndiffusion >>
rect 6 11 8 15
rect 10 11 12 15
rect 24 11 26 15
rect 28 11 30 15
rect 34 11 36 15
rect 38 11 40 15
rect 52 11 54 15
rect 56 11 64 15
rect 66 11 68 15
rect 80 11 82 15
rect 84 11 86 15
rect 90 11 92 15
rect 94 11 96 15
<< pdiffusion >>
rect 6 34 8 42
rect 10 34 12 42
rect 24 34 26 42
rect 28 34 36 42
rect 38 34 40 42
rect 52 34 54 42
rect 56 34 58 42
rect 62 34 64 42
rect 66 34 68 42
rect 80 34 82 42
rect 84 34 92 42
rect 94 34 96 42
<< metal1 >>
rect 0 52 102 53
rect 0 48 2 52
rect 6 48 20 52
rect 24 48 48 52
rect 52 48 68 52
rect 72 48 76 52
rect 80 48 102 52
rect 0 47 102 48
rect 2 42 6 47
rect 20 42 24 47
rect 48 42 52 47
rect 68 42 72 47
rect 76 42 80 47
rect 12 23 16 34
rect 40 23 44 34
rect 12 19 22 23
rect 30 19 50 23
rect 58 21 62 34
rect 96 30 100 34
rect 86 28 100 30
rect 70 26 100 28
rect 70 24 90 26
rect 12 15 16 19
rect 30 15 34 19
rect 58 17 72 21
rect 68 15 72 17
rect 86 15 90 24
rect 2 6 6 11
rect 20 6 24 11
rect 40 6 44 11
rect 48 6 52 11
rect 68 6 72 11
rect 76 6 80 11
rect 96 6 100 11
rect 0 5 103 6
rect 0 1 2 5
rect 6 1 20 5
rect 24 1 40 5
rect 44 1 48 5
rect 52 1 68 5
rect 72 1 76 5
rect 80 1 96 5
rect 100 1 103 5
rect 0 0 103 1
<< ntransistor >>
rect 8 11 10 15
rect 26 11 28 15
rect 36 11 38 15
rect 54 11 56 15
rect 64 11 66 15
rect 82 11 84 15
rect 92 11 94 15
<< ptransistor >>
rect 8 34 10 42
rect 26 34 28 42
rect 36 34 38 42
rect 54 34 56 42
rect 64 34 66 42
rect 82 34 84 42
rect 92 34 94 42
<< polycontact >>
rect 1 56 5 60
rect 22 19 26 23
rect 50 19 54 23
rect 66 24 70 28
rect 35 -7 39 -3
rect 81 -7 85 -3
<< ndcontact >>
rect 2 11 6 15
rect 12 11 16 15
rect 20 11 24 15
rect 30 11 34 15
rect 40 11 44 15
rect 48 11 52 15
rect 68 11 72 15
rect 76 11 80 15
rect 86 11 90 15
rect 96 11 100 15
rect 2 1 6 5
rect 20 1 24 5
rect 40 1 44 5
rect 48 1 52 5
rect 68 1 72 5
rect 76 1 80 5
rect 96 1 100 5
<< pdcontact >>
rect 2 48 6 52
rect 20 48 24 52
rect 48 48 52 52
rect 68 48 72 52
rect 76 48 80 52
rect 2 34 6 42
rect 12 34 16 42
rect 20 34 24 42
rect 40 34 44 42
rect 48 34 52 42
rect 58 34 62 42
rect 68 34 72 42
rect 76 34 80 42
rect 96 34 100 42
<< labels >>
rlabel metal1 32 52 32 52 1 VDD
rlabel metal1 60 3 60 3 1 GND
rlabel polycontact 37 -5 37 -5 1 Vin0
rlabel polycontact 83 -5 83 -5 1 Vin1
rlabel polycontact 3 58 3 58 3 Vselk
rlabel polysilicon 93 22 93 22 1 VselK
rlabel polycontact 24 21 24 21 1 snot
rlabel polycontact 52 21 52 21 1 and1
rlabel polycontact 68 26 68 26 1 and2
rlabel metal1 70 19 70 19 1 Vout
<< end >>
