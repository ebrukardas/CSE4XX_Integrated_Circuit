* SPICE3 file created from nor_8.ext - technology: scmos

.option scale=0.12u

M1000 a_n34_n18# VinA VDD w_n44_n24# pmos w=8 l=2
+  ad=64 pd=32 as=64 ps=44
M1001 Vout VinB a_n34_n18# w_n44_n24# pmos w=8 l=2
+  ad=48 pd=28 as=0 ps=0
M1002 Vout VinA GND Gnd nmos w=4 l=2
+  ad=32 pd=24 as=80 ps=72
M1003 GND VinB Vout Gnd nmos w=4 l=2
+  ad=0 pd=0 as=0 ps=0
C0 VinB w_n44_n24# 2.6fF
C1 VinA w_n44_n24# 2.6fF
C2 VDD w_n44_n24# 4.5fF
C3 Vout VinB 0.2fF
C4 Vout w_n44_n24# 1.9fF
C5 Vout Gnd 3.2fF
C6 VinB Gnd 5.6fF
C7 VinA Gnd 5.6fF
C8 VDD Gnd 3.6fF


*
* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    Vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2   V2   T3   V3   T4    V4    T5   V5    T5   V5     T5   V5     T5   V5 
*----- ----- ----- ------ --  --   ---  --   ---- --   ---   --    ---- --    ----  --    ----  --    ----  -- 
VinA   VinA   0    PWL(    0  0    3.9N  0   4N  2.5   7.9N  2.5   8N   0     11.9N  0     12N  2.5   15.9N  2.5  ) 
VinB   VinB   0    PWL(    0  0    3.9N  0   4N  0	   7.9N  0     8N   2.5   11.9N  2.5   12N  2.5   15.9N  2.5 )

*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  20.2N


* The following line is for DC analysis

.DC VINa 0 2.6 0.1

* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
