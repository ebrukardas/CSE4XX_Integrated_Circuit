* SPICE3 file created from inverter_8.ext - technology: scmos

.option scale=0.12u

M1000 Vout Vin VDD Vdd pmos w=8 l=2
+  ad=48 pd=28 as=64 ps=44
M1001 Vout Vin GND Gnd nmos w=4 l=2
+  ad=24 pd=20 as=40 ps=36
C0 Vdd Vin 2.6fF
C1 Vout Vdd 1.1fF
C2 Vdd VDD 3.7fF
C3 Vout Gnd 2.4fF
C4 Vin Gnd 5.6fF
C5 VDD Gnd 2.7fF


*
* INDEPENDANT VOLTAGE SOURCE
*
*Vname +NODE -NODE VALUE
*----- ----- ----- -----
VCC    Vdd     0     DC=2.5


* The following two lines are for TRANSIENT analysis
*
*Vname +Node -Node Option T1  V1   T2  V2   T3   V3   T4  V4  T5   V5 
*----- ----- ----- ------ --  --   --  --   ---- --   --  --  ---- -- 
Vin     Vin     0    PWL( 0   0    3.9N 0   4N   2.5  8N 2.5   8.1N  0  ) 



*     TSTEP TSTOP
*     ----- -----
.TRAN 0.1N  12N


* The following line is for DC analysis

.DC VIN 0 2.6 0.1

* TEMPERATURE and OPTIONS SETTING

.OPTIONS TEMP=25 reltol = 1e-6 

*MODELS

.include tsmc_cmos025

.END
